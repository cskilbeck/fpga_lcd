//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Wed Feb 14 11:53:37 2024

module Gowin_SP_text (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [11:0] ad;
input [7:0] din;

wire [27:0] sp_inst_0_dout_w;
wire [27:0] sp_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 4;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h00000003A407FCC56084970C48792705654302F60E904525F005618035452924;
defparam sp_inst_0.INIT_RAM_01 = 256'hE2359E570F941220104E1024E575C207E9431341F22010310D9807E9252D5D52;
defparam sp_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_03 = 256'h0000003720F94120EF0CC1205FA02F60E907E9CC960390F870CE1D018309B39E;
defparam sp_inst_0.INIT_RAM_04 = 256'h000000000000E2910EF0321540F40456FD03170CB5570398407F8304316B1522;
defparam sp_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_06 = 256'h0000004905EF4056180904E109230F407E9F7047E3170906C539D0F404913092;
defparam sp_inst_0.INIT_RAM_07 = 256'h00000000E325E5439C0DF2603571335D045F04152058303104913058302C53EF;
defparam sp_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_09 = 256'h000052FD02F6020F941204E1010F941203220EF037F8304543F80F870C487927;
defparam sp_inst_0.INIT_RAM_0A = 256'h000000000000E9606F05710584041091435540EF045940C3541354025F60E184;
defparam sp_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0C = 256'h005DD127F200914F403740F941204CF4095C9870FA055715CCF3020F94120398;
defparam sp_inst_0.INIT_RAM_0D = 256'h000000000000000E246123039806F025431D010317058204184091435E4570EF;
defparam sp_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_0F = 256'h325E5439C03EF9CC9D0F404E592604FF7DC55604E104E1970F94120A9215492F;
defparam sp_inst_0.INIT_RAM_10 = 256'h254E53520020F94120A4079C4E592604E10D217706F03592FD5D029584052183;
defparam sp_inst_0.INIT_RAM_11 = 256'h000F94120F40569C05CF8703980454F654058209604571035940487927056543;
defparam sp_inst_0.INIT_RAM_12 = 256'h000000E4913058302C9001805C0F5007E9B1D0317045F210452130580CC104E1;
defparam sp_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h0000EF024E575C207E9431341F2205840F407F83054529240104543F8095C987;
defparam sp_inst_0.INIT_RAM_15 = 256'h520F40257E124309256204C560490491304E107E9E565091435540EF020F9412;
defparam sp_inst_0.INIT_RAM_16 = 256'h0000000000000E2F710391409CEF204879270E553041805830E569704907E9F4;
defparam sp_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_18 = 256'h00045F2107E9BC1405418090C4130925604C5604E10321540E90CC1052570572;
defparam sp_inst_0.INIT_RAM_19 = 256'h00000000E5DD127F200914F405840EF04913058302C53E540431005840E90D98;
defparam sp_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1B = 256'h0041840914F404CF40CC520D1309B39E0254E53520010F9412025D2F607FCC56;
defparam sp_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000E2F94543010E90520F40E2F2031720487927;
defparam sp_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_1E = 256'h00000000003170418404E10C29105840EF03170580E58704521F304215803982;
defparam sp_inst_0.INIT_RAM_1F = 256'h00000000000000000000000000000000000000000000000000002E35F9714EF3;
defparam sp_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_21 = 256'h000000571D9088910E9045254390035BFF220FE52204E10415205B9D0C487927;
defparam sp_inst_0.INIT_RAM_22 = 256'h000000FE52204E10415205B9D0C4879270CEF940130571D901945D010C5325F3;
defparam sp_inst_0.INIT_RAM_23 = 256'h00007527043F804316B1522010F941204E52253088910E9045254390035BFF22;
defparam sp_inst_0.INIT_RAM_24 = 256'h04E104879270F4054529240108497091435E4570EF07F830398045E50F035D1A;
defparam sp_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000E235C7E9A06F07E9B205840310D980452923354;
defparam sp_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_27 = 256'h580ED98084970665430F9412045F21045F0425E04C5F30909B35C0F304C56092;
defparam sp_inst_0.INIT_RAM_28 = 256'h0039041840C3215900402F607E9A1D1031704E1030905840E907F83039840494;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000002ED9802F6056FC06F07E925F045F0E1083530390525840987;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h058408497048792704E104152045CC1307F830104543F8DF30F870C415205B9D;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000032204CF40C10F94120F40456FD09584052F6520F94120C13FC0EF0A4;
defparam sp_inst_0.INIT_RAM_2D = 256'h004104FF7204E10225431D7E92201031705804184091435E4570EF04316B1522;
defparam sp_inst_0.INIT_RAM_2E = 256'h000000000000000000000000000000000000000000000E2E905C0F5007E9CC50;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0F87094F25DF30435A04FE0E1D0F94120103170580C9C335C5294045B2F70582;
defparam sp_inst_0.INIT_RAM_31 = 256'h000000C4E9D03980E903170490E5DF804E5704E107F83058404940C05045E254;
defparam sp_inst_0.INIT_RAM_32 = 256'h00000000000000000000000000000000000000E23154906F07E9BE98403917C1;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h010F941205840DF26095C9D095C9D30310325E5439C0F40E7FEB0C35C9D09EF4;
defparam sp_inst_0.INIT_RAM_35 = 256'h001048792707E9CC130C4316B152203220EF0545292403980454410C7F8341F2;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000E2359E570F94122;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h000010EF0D98055304E105DF304C5F705C0F5006F034E135F8406F034524E582;
defparam sp_inst_0.INIT_RAM_39 = 256'h39807E97E92204E107E94139E5DDF306F09170398404180435A0580C7F8341F2;
defparam sp_inst_0.INIT_RAM_3A = 256'h00000000000000000000000000000000000E491305802C569C0F403254312183;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h000C48792705654304E109465C80359614092170395B3FA03394010F94120322;
defparam sp_inst_0.INIT_RAM_3D = 256'h0359614092170CEF940130571D903571D9094457C5325F30571D9048910C9201;
defparam sp_inst_0.INIT_RAM_3E = 256'h0004316B1522010F9412D85025E9830F42034355703980454E17048792704913;
defparam sp_inst_0.INIT_RAM_3F = 256'h00007E949270CD127143E90EF0545292401045218303E165039283043F807F83;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b00;
defparam sp_inst_1.BIT_WIDTH = 4;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h2222222744276666626767227666752676752766266266776726766276776675;
defparam sp_inst_1.INIT_RAM_01 = 256'h2277666626666722626662266666622666776666676262762666266676666667;
defparam sp_inst_1.INIT_RAM_02 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_03 = 256'h2222227232666652662666426652766266266666662762667226667664266664;
defparam sp_inst_1.INIT_RAM_04 = 256'h2222222222222766266277667267266766276722666727667276672776666676;
defparam sp_inst_1.INIT_RAM_05 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_06 = 256'h2222227626666267662426662776267266666272676724266677626726667242;
defparam sp_inst_1.INIT_RAM_07 = 256'h2222222227766677662667627666776627762666726672762666726672226666;
defparam sp_inst_1.INIT_RAM_08 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_09 = 256'h2222676627662326666526662326666524442662776672667766266722766675;
defparam sp_inst_1.INIT_RAM_0A = 256'h2222222222222332662666266727627667675266266662276666662776626667;
defparam sp_inst_1.INIT_RAM_0B = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_0C = 256'h2266667667727666527232666652666727666652642676666666232666652764;
defparam sp_inst_1.INIT_RAM_0D = 256'h2222222222222222276676276626627677662627672662276672766766665266;
defparam sp_inst_1.INIT_RAM_0E = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_0F = 256'h7766677642766666662672666676266662666626662766662666652377677664;
defparam sp_inst_1.INIT_RAM_10 = 256'h7676676772326666524422766666762666267672266276676666276667267667;
defparam sp_inst_1.INIT_RAM_11 = 256'h2226666726726666266667276626676766264223326666276662766675267675;
defparam sp_inst_1.INIT_RAM_12 = 256'h2222222666726672227776626676672666666276727766626676626626662666;
defparam sp_inst_1.INIT_RAM_13 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_14 = 256'h2222662266666622666776666676266726727667267766772626677662766665;
defparam sp_inst_1.INIT_RAM_15 = 256'h6626722666677727767227666276266672666266666762766767526623266665;
defparam sp_inst_1.INIT_RAM_16 = 256'h2222222222222226662776627666227666752666726662667266766276266666;
defparam sp_inst_1.INIT_RAM_17 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_18 = 256'h2227766626666667267662422667277672766626662776672662666267672652;
defparam sp_inst_1.INIT_RAM_19 = 256'h2222222226666766772766652667266266672667222676672776726672662666;
defparam sp_inst_1.INIT_RAM_1A = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_1B = 256'h2276672766652666726666766427666427676676772326666527667662766664;
defparam sp_inst_1.INIT_RAM_1C = 256'h2222222222222222222222222222226667772626626626726766276722766675;
defparam sp_inst_1.INIT_RAM_1D = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_1E = 256'h2222222222767276672666227662667266276726626667266766727766627642;
defparam sp_inst_1.INIT_RAM_1F = 256'h2222222222222222222222222222222222222222222222222222227766667666;
defparam sp_inst_1.INIT_RAM_20 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_21 = 256'h2222224444423333266266777667276666742667742666266652666422766675;
defparam sp_inst_1.INIT_RAM_22 = 256'h2222226677426662666526664227666752266677662666642444442452445545;
defparam sp_inst_1.INIT_RAM_23 = 256'h2222667427766277666667623266665276677742333326626677766727666674;
defparam sp_inst_1.INIT_RAM_24 = 256'h2666276667526726776677262676727667666652662766727662666676276664;
defparam sp_inst_1.INIT_RAM_25 = 256'h2222222222222222222222222227666666266266662266727626662666676766;
defparam sp_inst_1.INIT_RAM_26 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_27 = 256'h6422666267672667772666672776662776267662667662427667626727666242;
defparam sp_inst_1.INIT_RAM_28 = 256'h2276276672277667233276626667666276726662733266726627667276672666;
defparam sp_inst_1.INIT_RAM_29 = 256'h2222222222222222266627662676626626667767776266266772762676672767;
defparam sp_inst_1.INIT_RAM_2A = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_2B = 256'h2667267672766675266626665266666627667262667766266266722666526664;
defparam sp_inst_1.INIT_RAM_2C = 256'h2222222244426667223266665267266766276672676666266667266666266244;
defparam sp_inst_1.INIT_RAM_2D = 256'h2276266662266622767766666722627672662766727667666652662776666674;
defparam sp_inst_1.INIT_RAM_2E = 256'h2222222222222222222222222222222222222222222222266266766726666677;
defparam sp_inst_1.INIT_RAM_2F = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_30 = 256'h2667276666667277762766266626666726276726622767766676726667672642;
defparam sp_inst_1.INIT_RAM_31 = 256'h2222222666627662662767274226666276672666276672667266622772666777;
defparam sp_inst_1.INIT_RAM_32 = 256'h2222222222222222222222222222222222222222766662662666666672776766;
defparam sp_inst_1.INIT_RAM_33 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_34 = 256'h2326666526672667627666427666652762776667766267267666227666427665;
defparam sp_inst_1.INIT_RAM_35 = 256'h2262766675266666662277666667424442662677667727662666662276676667;
defparam sp_inst_1.INIT_RAM_36 = 256'h2222222222222222222222222222222222222222222222222227766662666672;
defparam sp_inst_1.INIT_RAM_37 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_38 = 256'h2222626626662667266626666266767266766726627666776672662766766742;
defparam sp_inst_1.INIT_RAM_39 = 256'h7662666666762666266676666766662662767276672666277762662276676667;
defparam sp_inst_1.INIT_RAM_3A = 256'h2222222222222222222222222222222222226667266222666626727767667666;
defparam sp_inst_1.INIT_RAM_3B = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam sp_inst_1.INIT_RAM_3C = 256'h2222766675267675266622766622766764277642776666626766232666652444;
defparam sp_inst_1.INIT_RAM_3D = 256'h2766764277642266677662666642544444255544244554524444423333266774;
defparam sp_inst_1.INIT_RAM_3E = 256'h2227766666762326666527422666672672277767627662667667276667526667;
defparam sp_inst_1.INIT_RAM_3F = 256'h2222666767722667667764266267766772626676672766742767642776627667;

endmodule //Gowin_SP_text
