//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Wed Feb 14 10:50:05 2024

module Gowin_SP_font (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [9:0] ad;
input [7:0] din;

wire [23:0] sp_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({gw_gnd,ad[9:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h0036367F367F3636000000000000363600180018183C3C180000000000000000;
defparam sp_inst_0.INIT_RAM_01 = 256'h0000000000030606006E333B6E1C361C0063660C18336300000C1F301E033E0C;
defparam sp_inst_0.INIT_RAM_02 = 256'h00000C0C3F0C0C000000663CFF3C660000060C1818180C0600180C0606060C18;
defparam sp_inst_0.INIT_RAM_03 = 256'h000103060C183060000C0C0000000000000000003F000000060C0C0000000000;
defparam sp_inst_0.INIT_RAM_04 = 256'h001E33301C30331E003F33061C30331E003F0C0C0C0C0E0C003E676F7B73633E;
defparam sp_inst_0.INIT_RAM_05 = 256'h000C0C0C1830333F001E33331F03061C001E3330301F033F0078307F33363C38;
defparam sp_inst_0.INIT_RAM_06 = 256'h060C0C00000C0C00000C0C00000C0C00000E18303E33331E001E33331E33331E;
defparam sp_inst_0.INIT_RAM_07 = 256'h000C000C1830331E00060C1830180C0600003F00003F000000180C0603060C18;
defparam sp_inst_0.INIT_RAM_08 = 256'h003C66030303663C003F66663E66663F0033333F33331E0C001E037B7B7B633E;
defparam sp_inst_0.INIT_RAM_09 = 256'h007C66730303663C000F06161E16467F007F46161E16467F001F36666666361F;
defparam sp_inst_0.INIT_RAM_0A = 256'h006766361E366667001E333330303078001E0C0C0C0C0C1E003333333F333333;
defparam sp_inst_0.INIT_RAM_0B = 256'h001C36636363361C006363737B6F67630063636B7F7F7763007F66460606060F;
defparam sp_inst_0.INIT_RAM_0C = 256'h001E33380E07331E006766363E66663F00381E3B3333331E000F06063E66663F;
defparam sp_inst_0.INIT_RAM_0D = 256'h0063777F6B636363000C1E3333333333003F333333333333001E0C0C0C0C2D3F;
defparam sp_inst_0.INIT_RAM_0E = 256'h001E06060606061E007F664C1831637F001E0C0C1E3333330063361C1C366363;
defparam sp_inst_0.INIT_RAM_0F = 256'hFF000000000000000000000063361C08001E18181818181E00406030180C0603;
defparam sp_inst_0.INIT_RAM_10 = 256'h001E3303331E0000003B66663E060607006E333E301E00000000000000180C0C;
defparam sp_inst_0.INIT_RAM_11 = 256'h1F303E33336E0000000F06060F06361C001E033F331E0000006E33333E303038;
defparam sp_inst_0.INIT_RAM_12 = 256'h0067361E366606071E33333030300030001E0C0C0C0E000C006766666E360607;
defparam sp_inst_0.INIT_RAM_13 = 256'h001E3333331E000000333333331F000000636B7F7F330000001E0C0C0C0C0C0E;
defparam sp_inst_0.INIT_RAM_14 = 256'h001F301E033E0000000F06666E3B000078303E33336E00000F063E66663B0000;
defparam sp_inst_0.INIT_RAM_15 = 256'h00367F7F6B630000000C1E3333330000006E33333333000000182C0C0C3E0C08;
defparam sp_inst_0.INIT_RAM_16 = 256'h00380C0C070C0C38003F260C193F00001F303E33333300000063361C36630000;
defparam sp_inst_0.INIT_RAM_17 = 256'h00000000000000000000000000003B6E00070C0C380C0C070018181800181818;

endmodule //Gowin_SP_font
